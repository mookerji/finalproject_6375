import Vector::*;
import TomasuloTypes::*;
import FShow::*;
import ReorderBuffer::*;

interface ReservationStation;
  method ActionValue#(RSEntry) getReadyEntry();
  method Action put(RSEntry entry);
endinterface

module mkReservationStation(ROB#(16) rob, ReservationStation rsifc);

  Vector#(2, Reg#(Maybe#(RSEntry))) entries <- replicateM(mkReg(tagged Invalid));

/*
  rule fucklife;
    for (Integer i = 0; i < 2; i = i + 1) begin
      case (entries[i]) matches
        tagged Valid .e: $display("Reservation Station contains entry ",fshow(e.op)," [",fshow(e.op1),", ",fshow(e.op2),"]");
        tagged Invalid: $display("Reservation Station contains no entry");
      endcase
    end
  endrule
*/

  rule allfull(isValid(entries[0]) && isValid(entries[1]));
    $display("oscar the grouch lives in a trashcan");
  endrule

  rule check_for_completion_of_dependencies;
$display("RS Check start");
    for (Integer i = 0; i < 2; i = i + 1) begin
      if (isValid(entries[i])) begin
        let entry = fromMaybe(?, entries[i]);
        Bool modified = False;
$display("Looking for ",fshow(entry.op1));
if (entry.op1 matches tagged Tag .it) $display("data for the above tag in the ROB is ",rob.get(it));
        if (entry.op1 matches tagged Tag .it &&& rob.get(it) matches tagged Valid .robent &&&
            robent.data matches tagged Valid .robdata) begin
           entry.op1 = tagged Imm robdata;
           modified = True;
        end
$display("Looking for ",fshow(entry.op2));
if (entry.op2 matches tagged Tag .it) $display("data for the above tag in the ROB is ",rob.get(it));
        if (entry.op2 matches tagged Tag .it &&& rob.get(it) matches tagged Valid .robent &&&
            robent.data matches tagged Valid .robdata) begin
           entry.op2 = tagged Imm robdata;
           modified = True;
        end
        if (modified) begin
          $display("Reservation Station found ROB update which updated an RSEntry");
          entries[i] <= tagged Valid entry;
        end
      end
    end
$display("RS Check end");
  endrule

  function Maybe#(UInt#(TLog#(2))) readyEntry();
    Maybe#(UInt#(TLog#(2))) index = tagged Invalid;
    for (Integer i = 0; i < 2; i = i + 1) begin
      if (isValid(entries[i])) begin
        let entry = fromMaybe(?, entries[i]);
        if (entry.op1 matches tagged Imm .a &&& entry.op2 matches tagged Imm .b) begin
          index = tagged Valid fromInteger(i);
        end
      end
    end
    return index;
  endfunction

  function Maybe#(UInt#(TLog#(2))) freeSlot();
    Maybe#(UInt#(TLog#(2))) index = tagged Invalid;
    for (Integer i = 0; i < 2; i = i + 1) begin
      if (!isValid(entries[i])) begin
        index = tagged Valid fromInteger(i);
      end
    end
    return index;
  endfunction

  method ActionValue#(RSEntry) getReadyEntry() if (readyEntry() matches tagged Valid .i);
    let e = fromMaybe(?, entries[i]);
    entries[i] <= tagged Invalid;
    $display("Got ready entry ",fshow(e.op)," [",fshow(e.op1),", ",fshow(e.op2),"]");
    return e;
  endmethod

  method Action put(RSEntry entry) if (isValid(freeSlot()));
    let i = fromMaybe(?, readyEntry());
    entries[i] <= tagged Valid entry;
  endmethod
endmodule
